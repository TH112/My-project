
module system (
	clk_clk,
	hex_0_conduit_end_hex,
	reset_reset_n,
	switch_0_conduit_end_export);	

	input		clk_clk;
	output	[6:0]	hex_0_conduit_end_hex;
	input		reset_reset_n;
	input	[31:0]	switch_0_conduit_end_export;
endmodule
